// Code your testbench here
// or browse Examples
module testbench();
  logic clk;
  logic reset;
  logic [31:0] WriteData, DataAdr;
  logic MemWrite;    // instantiate device to be tested    
  
  top dut(clk, reset, WriteData, DataAdr, MemWrite);    // initialize test    
  
  initial      
    begin           
      reset <= 1; # 22; reset <= 0;
    end    // generate clock to sequence tests    
	 
  always    
    begin           
    clk <= 1; # 5; clk <= 0; # 5;    
    end    // check results    
	 
  always @(negedge clk)   
    begin           
      if(MemWrite) 
        begin
        if(DataAdr === 100 & WriteData === 25) 
          begin              $display("Simulation succeeded");
            $stop;
          end 
          else if (DataAdr !== 96)
            begin              
              $display("Simulation failed");
              $stop;
            end
        end
      end
endmodule



module top(input   logic clk, reset,
           output logic [31:0] WriteData, DataAdr,
           output logic             MemWrite);
  logic [31:0] PC, Instr, ReadData;    // instantiate processor and memories      
  riscvsingle rvsingle( clk, reset, PC, Instr, MemWrite, DataAdr,  WriteData, ReadData);
  imem imem(PC, Instr);    
  dmem dmem(clk, MemWrite, DataAdr, WriteData, ReadData);
endmodule

module imem(input     logic [31:0] a,
            output logic [31:0] rd);
  logic [31:0] RAM[63:0];
  assign RAM[0] = 32'h00500113;
  assign RAM[1] = 32'h00C00193;
  initial       
	begin
	$readmemh("riscvtest.txt",RAM);
	//assign RAM[0] = 32'h00500113;
	end
  assign rd = RAM[a[31:2]];
  // word aligned
endmodule

module dmem(input     logic clk, we,
            input     logic [31:0] a, wd,
            output logic [31:0] rd);
  logic [31:0] RAM[63:0];
  
  assign rd = RAM[a[31:2]]; // word aligned    

  always_ff @(posedge clk)
    if (we) RAM[a[31:2]] <= wd;
endmodule

