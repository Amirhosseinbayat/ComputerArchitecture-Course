module ControlBufferRegister();

endmodule
