module SequentialLogic();

endmodule
