module ControlMemory();

endmodule
